module ForwardSbox(
	input [7:0] data,
	output reg [7:0] fsb_data
);

always@(*) begin
	case(data)
		// data[7:4] = 4'h0
		8'h00: fsb_data = 8'h63;
		8'h01: fsb_data = 8'h7c;
		8'h02: fsb_data = 8'h77;
		8'h03: fsb_data = 8'h7b;
		8'h04: fsb_data = 8'hf2;
		8'h05: fsb_data = 8'h6b;
		8'h06: fsb_data = 8'h6f;
		8'h07: fsb_data = 8'hc5;
		8'h08: fsb_data = 8'h30;
		8'h09: fsb_data = 8'h01;
		8'h0a: fsb_data = 8'h67;
		8'h0b: fsb_data = 8'h2b;
		8'h0c: fsb_data = 8'hfe;
		8'h0d: fsb_data = 8'hd7;
		8'h0e: fsb_data = 8'hab;
		8'h0f: fsb_data = 8'h76;
		// data[7:4] = 4'h1
		8'h10: fsb_data = 8'hca;
		8'h11: fsb_data = 8'h82;
		8'h12: fsb_data = 8'hc9;
		8'h13: fsb_data = 8'h7d;
		8'h14: fsb_data = 8'hfa;
		8'h15: fsb_data = 8'h59;
		8'h16: fsb_data = 8'h47;
		8'h17: fsb_data = 8'hf0;
		8'h18: fsb_data = 8'had;
		8'h19: fsb_data = 8'hd4;
		8'h1a: fsb_data = 8'ha2;
		8'h1b: fsb_data = 8'haf;
		8'h1c: fsb_data = 8'h9c;
		8'h1d: fsb_data = 8'ha4;
		8'h1e: fsb_data = 8'h72;
		8'h1f: fsb_data = 8'hc0;
		// data[7:4] = 4'h2
		8'h20: fsb_data = 8'hb7;
		8'h21: fsb_data = 8'hfd;
		8'h22: fsb_data = 8'h93;
		8'h23: fsb_data = 8'h26;
		8'h24: fsb_data = 8'h36;
		8'h25: fsb_data = 8'h3f;
		8'h26: fsb_data = 8'hf7;
		8'h27: fsb_data = 8'hcc;
		8'h28: fsb_data = 8'h34;
		8'h29: fsb_data = 8'ha5;
		8'h2a: fsb_data = 8'he5;
		8'h2b: fsb_data = 8'hf1;
		8'h2c: fsb_data = 8'h71;
		8'h2d: fsb_data = 8'hd8;
		8'h2e: fsb_data = 8'h31;
		8'h2f: fsb_data = 8'h15;
		// data[7:4] = 4'h3
		8'h30: fsb_data = 8'h04;
		8'h31: fsb_data = 8'hc7;
		8'h32: fsb_data = 8'h23;
		8'h33: fsb_data = 8'hc3;
		8'h34: fsb_data = 8'h18;
		8'h35: fsb_data = 8'h96;
		8'h36: fsb_data = 8'h05;
		8'h37: fsb_data = 8'h9a;
		8'h38: fsb_data = 8'h07;
		8'h39: fsb_data = 8'h12;
		8'h3a: fsb_data = 8'h80;
		8'h3b: fsb_data = 8'he2;
		8'h3c: fsb_data = 8'heb;
		8'h3d: fsb_data = 8'h27;
		8'h3e: fsb_data = 8'hb2;
		8'h3f: fsb_data = 8'h75;
		// data[7:4] = 4'h4
		8'h40: fsb_data = 8'h09;
		8'h41: fsb_data = 8'h83;
		8'h42: fsb_data = 8'h2c;
		8'h43: fsb_data = 8'h1a;
		8'h44: fsb_data = 8'h1b;
		8'h45: fsb_data = 8'h6e;
		8'h46: fsb_data = 8'h5a;
		8'h47: fsb_data = 8'ha0;
		8'h48: fsb_data = 8'h52;
		8'h49: fsb_data = 8'h3b;
		8'h4a: fsb_data = 8'hd6;
		8'h4b: fsb_data = 8'hb3;
		8'h4c: fsb_data = 8'h29;
		8'h4d: fsb_data = 8'he3;
		8'h4e: fsb_data = 8'h2f;
		8'h4f: fsb_data = 8'h84;
		// data[7:4] = 4'h5
		8'h50: fsb_data = 8'h53;
		8'h51: fsb_data = 8'hd1;
		8'h52: fsb_data = 8'h00;
		8'h53: fsb_data = 8'hed;
		8'h54: fsb_data = 8'h20;
		8'h55: fsb_data = 8'hfc;
		8'h56: fsb_data = 8'hb1;
		8'h57: fsb_data = 8'h5b;
		8'h58: fsb_data = 8'h6a;
		8'h59: fsb_data = 8'hcb;
		8'h5a: fsb_data = 8'hbe;
		8'h5b: fsb_data = 8'h39;
		8'h5c: fsb_data = 8'h4a;
		8'h5d: fsb_data = 8'h4c;
		8'h5e: fsb_data = 8'h58;
		8'h5f: fsb_data = 8'hcf;
		// data[7:4] = 4'h6
		8'h60: fsb_data = 8'hd0;
		8'h61: fsb_data = 8'hef;
		8'h62: fsb_data = 8'haa;
		8'h63: fsb_data = 8'hfb;
		8'h64: fsb_data = 8'h43;
		8'h65: fsb_data = 8'h4d;
		8'h66: fsb_data = 8'h33;
		8'h67: fsb_data = 8'h85;
		8'h68: fsb_data = 8'h45;
		8'h69: fsb_data = 8'hf9;
		8'h6a: fsb_data = 8'h02;
		8'h6b: fsb_data = 8'h7f;
		8'h6c: fsb_data = 8'h50;
		8'h6d: fsb_data = 8'h3c;
		8'h6e: fsb_data = 8'h9f;
		8'h6f: fsb_data = 8'ha8;
		// data[7:4] = 4'h7
		8'h70: fsb_data = 8'h51;
		8'h71: fsb_data = 8'ha3;
		8'h72: fsb_data = 8'h40;
		8'h73: fsb_data = 8'h8f;
		8'h74: fsb_data = 8'h92;
		8'h75: fsb_data = 8'h9d;
		8'h76: fsb_data = 8'h38;
		8'h77: fsb_data = 8'hf5;
		8'h78: fsb_data = 8'hbc;
		8'h79: fsb_data = 8'hb6;
		8'h7a: fsb_data = 8'hda;
		8'h7b: fsb_data = 8'h21;
		8'h7c: fsb_data = 8'h10;
		8'h7d: fsb_data = 8'hff;
		8'h7e: fsb_data = 8'hf3;
		8'h7f: fsb_data = 8'hd2;
		// data[7:4] = 4'h8
		8'h80: fsb_data = 8'hcd;
		8'h81: fsb_data = 8'h0c;
		8'h82: fsb_data = 8'h13;
		8'h83: fsb_data = 8'hec;
		8'h84: fsb_data = 8'h5f;
		8'h85: fsb_data = 8'h97;
		8'h86: fsb_data = 8'h44;
		8'h87: fsb_data = 8'h17;
		8'h88: fsb_data = 8'hc4;
		8'h89: fsb_data = 8'ha7;
		8'h8a: fsb_data = 8'h7e;
		8'h8b: fsb_data = 8'h3d;
		8'h8c: fsb_data = 8'h64;
		8'h8d: fsb_data = 8'h5d;
		8'h8e: fsb_data = 8'h19;
		8'h8f: fsb_data = 8'h73;
		// data[7:4] = 4'h9
		8'h90: fsb_data = 8'h60;
		8'h91: fsb_data = 8'h81;
		8'h92: fsb_data = 8'h4f;
		8'h93: fsb_data = 8'hdc;
		8'h94: fsb_data = 8'h22;
		8'h95: fsb_data = 8'h2a;
		8'h96: fsb_data = 8'h90;
		8'h97: fsb_data = 8'h88;
		8'h98: fsb_data = 8'h46;
		8'h99: fsb_data = 8'hee;
		8'h9a: fsb_data = 8'hb8;
		8'h9b: fsb_data = 8'h14;
		8'h9c: fsb_data = 8'hde;
		8'h9d: fsb_data = 8'h5e;
		8'h9e: fsb_data = 8'h0b;
		8'h9f: fsb_data = 8'hdb;
		// data[7:4] = 4'ha
		8'ha0: fsb_data = 8'he0;
		8'ha1: fsb_data = 8'h32;
		8'ha2: fsb_data = 8'h3a;
		8'ha3: fsb_data = 8'h0a;
		8'ha4: fsb_data = 8'h49;
		8'ha5: fsb_data = 8'h06;
		8'ha6: fsb_data = 8'h24;
		8'ha7: fsb_data = 8'h5c;
		8'ha8: fsb_data = 8'hc2;
		8'ha9: fsb_data = 8'hd3;
		8'haa: fsb_data = 8'hac;
		8'hab: fsb_data = 8'h62;
		8'hac: fsb_data = 8'h91;
		8'had: fsb_data = 8'h95;
		8'hae: fsb_data = 8'he4;
		8'haf: fsb_data = 8'h79;
		// data[7:4] = 4'hb
		8'hb0: fsb_data = 8'he7;
		8'hb1: fsb_data = 8'hc8;
		8'hb2: fsb_data = 8'h37;
		8'hb3: fsb_data = 8'h6d;
		8'hb4: fsb_data = 8'h8d;
		8'hb5: fsb_data = 8'hd5;
		8'hb6: fsb_data = 8'h4e;
		8'hb7: fsb_data = 8'ha9;
		8'hb8: fsb_data = 8'h6c;
		8'hb9: fsb_data = 8'h56;
		8'hba: fsb_data = 8'hf4;
		8'hbb: fsb_data = 8'hea;
		8'hbc: fsb_data = 8'h65;
		8'hbd: fsb_data = 8'h7a;
		8'hbe: fsb_data = 8'hae;
		8'hbf: fsb_data = 8'h08;
		// data[7:4] = 4'hc
		8'hc0: fsb_data = 8'hba;
		8'hc1: fsb_data = 8'h78;
		8'hc2: fsb_data = 8'h25;
		8'hc3: fsb_data = 8'h2e;
		8'hc4: fsb_data = 8'h1c;
		8'hc5: fsb_data = 8'ha6;
		8'hc6: fsb_data = 8'hb4;
		8'hc7: fsb_data = 8'hc6;
		8'hc8: fsb_data = 8'he8;
		8'hc9: fsb_data = 8'hdd;
		8'hca: fsb_data = 8'h74;
		8'hcb: fsb_data = 8'h1f;
		8'hcc: fsb_data = 8'h4b;
		8'hcd: fsb_data = 8'hbd;
		8'hce: fsb_data = 8'h8b;
		8'hcf: fsb_data = 8'h8a;
		// data[7:4] = 4'hd
		8'hd0: fsb_data = 8'h70;
		8'hd1: fsb_data = 8'h3e;
		8'hd2: fsb_data = 8'hb5;
		8'hd3: fsb_data = 8'h66;
		8'hd4: fsb_data = 8'h48;
		8'hd5: fsb_data = 8'h03;
		8'hd6: fsb_data = 8'hf6;
		8'hd7: fsb_data = 8'h0e;
		8'hd8: fsb_data = 8'h61;
		8'hd9: fsb_data = 8'h35;
		8'hda: fsb_data = 8'h57;
		8'hdb: fsb_data = 8'hb9;
		8'hdc: fsb_data = 8'h86;
		8'hdd: fsb_data = 8'hc1;
		8'hde: fsb_data = 8'h1d;
		8'hdf: fsb_data = 8'h9e;
		// data[7:4] = 4'he
		8'he0: fsb_data = 8'he1;
		8'he1: fsb_data = 8'hf8;
		8'he2: fsb_data = 8'h98;
		8'he3: fsb_data = 8'h11;
		8'he4: fsb_data = 8'h69;
		8'he5: fsb_data = 8'hd9;
		8'he6: fsb_data = 8'h8e;
		8'he7: fsb_data = 8'h94;
		8'he8: fsb_data = 8'h9b;
		8'he9: fsb_data = 8'h1e;
		8'hea: fsb_data = 8'h87;
		8'heb: fsb_data = 8'he9;
		8'hec: fsb_data = 8'hce;
		8'hed: fsb_data = 8'h55;
		8'hee: fsb_data = 8'h28;
		8'hef: fsb_data = 8'hdf;
		// data[7:4] = 4'hf
		8'hf0: fsb_data = 8'h8c;
		8'hf1: fsb_data = 8'ha1;
		8'hf2: fsb_data = 8'h89;
		8'hf3: fsb_data = 8'h0d;
		8'hf4: fsb_data = 8'hbf;
		8'hf5: fsb_data = 8'he6;
		8'hf6: fsb_data = 8'h42;
		8'hf7: fsb_data = 8'h68;
		8'hf8: fsb_data = 8'h41;
		8'hf9: fsb_data = 8'h99;
		8'hfa: fsb_data = 8'h2d;
		8'hfb: fsb_data = 8'h0f;
		8'hfc: fsb_data = 8'hb0;
		8'hfd: fsb_data = 8'h54;
		8'hfe: fsb_data = 8'hbb;
		8'hff: fsb_data = 8'h16;
	endcase
end

endmodule